/* @wavedrom 
{
    signal : [
        { name: "clk",  wave: "P....................", phase: 0, period: 1},
        { name: "rstn",  wave: "0.1..................", phase: 0, period: 1},
    ]
}
*/
`timescale 1ns/1ps

module tb_top;

//------------------------------------------
// �ź�����
//------------------------------------------
    reg        	    clk;
    reg [4:0]       Wr_idx;
    reg [4:0]       R1_idx;
    reg [4:0]       R2_idx;
    reg [31:0]      Data_in;
    reg             Wr_en;

    wire [31:0] 	REG_1;
    wire [31:0] 	REG_2;
//------------------------------------------
// ʵ����������ģ��
//------------------------------------------
top u_top(
	.clk     	( clk      ),
	.Wr_idx  	( Wr_idx   ),
	.R1_idx  	( R1_idx   ),
	.R2_idx  	( R2_idx   ),
	.Data_in 	( Data_in  ),
	.Wr_en   	( Wr_en    ),

	.REG_1   	( REG_1    ),
	.REG_2   	( REG_2    )
);

//------------------------------------------
// ����ʱ�ӣ�20ns, 50MHz
//------------------------------------------
    initial begin
        clk = 1;
        forever #10 clk = ~clk;
    end
//------------------------------------------
// ��λ
//------------------------------------------

//------------------------------------------
// Test sequence
//------------------------------------------

    initial begin
        $dumpfile("tb_top.vcd");
        $dumpvars(0, tb_top);

        #5;     // Wait for a few time units
        Wr_idx = 5'd1;   
        R1_idx = 5'd0;
        R2_idx = 5'd0;
        Data_in = 32'hDEAD_BEEF;
        Wr_en = 1;
        #20;
        Wr_idx = 5'd2;   
        R1_idx = 5'd0;
        R2_idx = 5'd0;
        Data_in = 32'h1234_5678;
        Wr_en = 1;
        #20;
        Wr_idx = 5'd0;   
        R1_idx = 5'd1;
        R2_idx = 5'd2;
        Data_in = 32'h0000_0000;
        Wr_en = 0;
        #20;

        #100;
        $finish;
    end
    
endmodule


