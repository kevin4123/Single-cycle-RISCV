`timescale 1ns/1ps

module tb_top;

//------------------------------------------
// �ź�����
//------------------------------------------
    reg [31:0]      Addr;

    wire [31:0] 	Instr;
//------------------------------------------
// ʵ����������ģ��
//------------------------------------------
top u_top(
	.Addr  	( Addr   ),
	.Instr 	( Instr  )
);
//------------------------------------------
// ����ʱ�ӣ�20ns, 50MHz
//------------------------------------------

//------------------------------------------
// ��λ
//------------------------------------------

//------------------------------------------
// Test sequence
//------------------------------------------

    initial begin
        $dumpfile("tb_top.vcd");
        $dumpvars(0, tb_top);

        #5;     // Wait for a few time units  
        Addr = 32'h0300_0000;   // outside cs: 0
        #20;
        Addr = 32'h0400_0000;   // 0
        #20;
        Addr = 32'h0400_0004;   // 1
        #20;
        Addr = 32'h0400_0008;   // 2
        #20;
        Addr = 32'h0400_0009;   // 2 (unaligned)

        #100;
        $finish;
    end
    
endmodule


